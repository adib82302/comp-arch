    Mac OS X            	   2   �      �                                      ATTR       �   �   (                  �     com.apple.lastuseddate#PS       �     com.apple.quarantine ���g    ��H1    q/0086;67a3acf6;BBEdit; 