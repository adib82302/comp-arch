    Mac OS X            	   2   �      �                                      ATTR       �   �   (                  �     com.apple.lastuseddate#PS       �     com.apple.quarantine 4ۤg    ��!    q/0086;67a4db34;BBEdit; 