// This file has the parameter and typedefs used in lab 3 part b

`ifndef __SYS_DEFS_VH__
`define __SYS_DEFS_VH__

typedef enum logic [1:0] {WAIT, WATCH, ASSERT} STATE;
typedef enum logic [1:0] {RAND, MATCH, NO_MATCH} OVERRIDE;

`endif // __SYS_DEFS_VH__
