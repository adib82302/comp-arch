    Mac OS X            	   2   �      �                                      ATTR       �   �   (                  �     com.apple.lastuseddate#PS       �     com.apple.quarantine 7ۤg    X��    q/0086;67a4db37;BBEdit; 